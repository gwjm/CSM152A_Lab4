`timescale 1ns/1ps


module SPIControl(
    clk,
    rst,
    sndRec,
    busy,
    dSend,
    RxData,
    ss,
    getByte,
    sndData,
    dread
);

endmodule