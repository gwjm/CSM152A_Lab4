`timescale 1ns/1ps

module PMODJSTK(
    clk, 
    rst, 
    sndrcv,
    dsend, 
    miso, 
    ss,
    sclk,
    mosi,
    dread
);

endmodule 