`timescale 1ns/1ps

module SPI_Interface(
    clk,
    rst,
    sndRec,
    dSend,
    miso,
    mosi,
    sclk,
	busy,
    dread
);

endmodule